////////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   / 
// /___/  \  /    Vendor: Xilinx 
// \   \   \/     Version : 3.5
//  \   \         Application : 7 Series FPGAs Transceivers Wizard 
//  /   /         Filename : gtwizard_0_rx_manual_phase_align.v
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\ 
//
//
//  Description :     This module performs RX Buffer Phase Alignment in Manual Mode.
//                     
//
//
// Module gtwizard_0_rx_manual_phase_align
// Generated by Xilinx 7 Series FPGAs Transceivers Wizard
// 
// 
// (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES. 



`timescale 1ns / 1ps
`define DLY #1

module gtwizard_0_RX_MANUAL_PHASE_ALIGN  #
  (
    parameter NUMBER_OF_LANES = 4,  // Number of lanes that are controlled using this FSM.
    parameter MASTER_LANE_ID  = 0   // Number of the lane which is considered the master 
                                    // in manual phase-alignment
   )
   (
    input   wire                             STABLE_CLOCK,              //Stable Clock, either a stable clock from the PCB
    input   wire                             RESET_PHALIGNMENT,
    input   wire                             RUN_PHALIGNMENT,
    output  reg                              PHASE_ALIGNMENT_DONE = 1'b0,      // Manual phase-alignment performed sucessfully    
    output  reg     [NUMBER_OF_LANES-1:0]    RXDLYSRESET = {NUMBER_OF_LANES{1'b0}},              
    input   wire    [NUMBER_OF_LANES-1:0]    RXDLYSRESETDONE,          
    output  reg     [NUMBER_OF_LANES-1:0]    RXPHALIGN = {NUMBER_OF_LANES{1'b0}},                
    input   wire    [NUMBER_OF_LANES-1:0]    RXPHALIGNDONE,
    output  reg     [NUMBER_OF_LANES-1:0]    RXDLYEN = {NUMBER_OF_LANES{1'b0}}                  
    );
              
           
   genvar j;
   integer i;
   wire [NUMBER_OF_LANES-1:0] VCC_VEC = {NUMBER_OF_LANES{1'b1}};
   wire [NUMBER_OF_LANES-1:0] GND_VEC = {NUMBER_OF_LANES{1'b0}};

   localparam [2:0]
               INIT             = 3'b000,
               WAIT_DLYRST_DONE = 3'b001,
               M_PHALIGN        = 3'b010,
               M_DLYEN          = 3'b011,
               S_PHALIGN        = 3'b100,
               M_DLYEN2         = 3'b101,
               PHALIGN_DONE     = 3'b110;

  reg [2:0] rx_phalign_manual_state = INIT;


  reg  [NUMBER_OF_LANES-1:0] rxphaligndone_prev = {NUMBER_OF_LANES{1'b0}};
  wire [NUMBER_OF_LANES-1:0] rxphaligndone_ris_edge;
  reg  [NUMBER_OF_LANES-1:0] rxdlysresetdone_store= {NUMBER_OF_LANES{1'b0}};
  reg  [NUMBER_OF_LANES-1:0] rxphaligndone_store = {NUMBER_OF_LANES{1'b0}};
  reg                        rxdone_clear = 1'b0;
  wire [NUMBER_OF_LANES-1:0] rxphaligndone_sync; 
  wire [NUMBER_OF_LANES-1:0] rxdlysresetdone_sync; 


  //Clock Domain Crossing

 generate
  for (j = 0;j <= NUMBER_OF_LANES-1;j = j+1) begin

 gtwizard_0_sync_block sync_RXPHALIGNDONE
        (
           .clk             (STABLE_CLOCK),
           .data_in         (RXPHALIGNDONE[j]),
           .data_out        (rxphaligndone_sync[j])
        );

 gtwizard_0_sync_block sync_RXDLYSRESETDONE
        (
           .clk             (STABLE_CLOCK),
           .data_in         (RXDLYSRESETDONE[j]),
           .data_out        (rxdlysresetdone_sync[j])
        );
  end 
 endgenerate

  always @(posedge STABLE_CLOCK)
  begin
      rxphaligndone_prev    <= `DLY  rxphaligndone_sync;  
  end 
 
 generate 
   for (j = 0;j <=  NUMBER_OF_LANES-1;j = j+1)
   begin
    assign  rxphaligndone_ris_edge[j] = ((rxphaligndone_prev[j] == 1'b0) && (rxphaligndone_sync[j] == 1'b1))  ? 1'b1 : 1'b0;            
   end
  endgenerate


  always @(posedge STABLE_CLOCK)
  begin
      if (rxdone_clear) 
      begin
        rxdlysresetdone_store <= `DLY  GND_VEC;
        rxphaligndone_store   <= `DLY  GND_VEC;
      end

      else
      begin
        for (i = 0; i <= NUMBER_OF_LANES-1; i = i+1) 
        begin
          if (rxdlysresetdone_sync[i] == 1'b1)
            rxdlysresetdone_store[i] <= `DLY  1'b1;

          if (rxphaligndone_ris_edge[i] == 1'b1)
             rxphaligndone_store[i]  <= `DLY  1'b1;
        end 
      end
  end




  always @(posedge STABLE_CLOCK)
  begin
      if (RESET_PHALIGNMENT == 1)
      begin
        PHASE_ALIGNMENT_DONE    <= `DLY  1'b0;
        RXDLYSRESET             <= `DLY  {NUMBER_OF_LANES{1'b0}};
        RXPHALIGN               <= `DLY  {NUMBER_OF_LANES{1'b0}};
        RXDLYEN                 <= `DLY  {NUMBER_OF_LANES{1'b0}};
        rx_phalign_manual_state <= `DLY  INIT;
        rxdone_clear            <= `DLY  1'b1;

      end
      else
      begin
        case (rx_phalign_manual_state)
           INIT :
           begin 
            PHASE_ALIGNMENT_DONE <= `DLY  1'b0;
            rxdone_clear         <= `DLY  1'b1;

            if (RUN_PHALIGNMENT)
            begin
              //Assert RXDLYSRESET for all lanes. 
              rxdone_clear            <= `DLY  1'b0;
              RXDLYSRESET             <= `DLY  {NUMBER_OF_LANES{1'b1}};
              rx_phalign_manual_state <= `DLY  WAIT_DLYRST_DONE;
            end
           end
            
           WAIT_DLYRST_DONE :
           begin
            for (i = 0;i <= NUMBER_OF_LANES - 1;i = i+1)
            begin
              if (rxdlysresetdone_store[i] == 1) 
                //Hold RXDLYSRESET High until RXDLYSRESETDONE of the 
                //respective lane is asserted.
                //Deassert RXDLYSRESET for the lane in which the 
                //RXDLYSRESETDONE is asserted.
                RXDLYSRESET[i] <= `DLY  0;
            end
            if (rxdlysresetdone_store == VCC_VEC)
            begin
              rx_phalign_manual_state   <= `DLY  M_PHALIGN;
            end
           end
          
           M_PHALIGN :
           begin 
            //When RXDLYSRESET of all lanes are deasserted, assert 
            //RXPHALIGN for the master lane.
            RXPHALIGN[MASTER_LANE_ID] <= `DLY  1'b1;
            if (rxphaligndone_ris_edge[MASTER_LANE_ID] == 1)
            begin
              //Hold this signal High until a rising edge on RXPHALIGNDONE 
              //of the master lane is detected, then deassert RXPHALIGN for 
              //the master lane.
              RXPHALIGN[MASTER_LANE_ID] <= `DLY  1'b0;
              rx_phalign_manual_state   <= `DLY  M_DLYEN;
            end
           end
          
           M_DLYEN :
           begin 
            //Assert RXDLYEN for the master lane. This causes RXPHALIGNDONE 
            //to be deasserted.
            RXDLYEN[MASTER_LANE_ID] <= `DLY  1'b1;
            if (rxphaligndone_ris_edge[MASTER_LANE_ID] == 1)
            begin
              //Hold RXDLYEN for the master lane High until a rising edge on
              //RXPHALIGNDONE of the master lane is detected, then deassert 
              //RXDLYEN for the master lane.
              RXDLYEN[MASTER_LANE_ID]   <= `DLY  1'b0;
              rx_phalign_manual_state   <= `DLY  S_PHALIGN;  
            end
           end
          
           S_PHALIGN :
           begin
            //Assert RXPHALIGN for all slave lane(s). Hold this signal High until
            //a rising edge on RXPHALIGNDONE of the respective slave lane is detected.
            RXPHALIGN                 <= `DLY  {NUMBER_OF_LANES{1'b1}};//\Assert only the PHINIT-signal of
            RXPHALIGN[MASTER_LANE_ID] <= `DLY  0;          ///the slaves.
            for (i = 0;i <=  NUMBER_OF_LANES - 1;i = i+1)
            begin
              if (rxphaligndone_store[i] == 1)
                //When a rising edge on the respective lane is detected, RXPHALIGN
                //of that lane is deasserted.
                RXPHALIGN[i] <= `DLY  1'b0;
            end 
           //The reason for checking of the occurance of at least one rising edge
            //is to avoid the potential direct move where RXPHALIGNDONE might not 
            //be going low fast enough. 
            if (rxphaligndone_store == VCC_VEC) 
              rx_phalign_manual_state   <= `DLY  M_DLYEN2;
           end
          
           M_DLYEN2 :
           begin
            //When RXPHALIGN for all slave lane(s) are deasserted, assert RXDLYEN 
            //for the master lane. This causes RXPHALIGNDONE of the master lane 
            //to be deasserted.
            RXDLYEN[MASTER_LANE_ID] <= `DLY  1'b1;
            if (rxphaligndone_ris_edge[MASTER_LANE_ID] == 1)
              //Wait until RXPHALIGNDONE of the master lane reasserts. Phase and 
              //delay alignment for the multilane interface is complete.
              rx_phalign_manual_state   <= `DLY  PHALIGN_DONE;        
           end 
          
           PHALIGN_DONE :
           begin
            //Continue to hold RXDLYEN for the master lane High to adjust RXUSRCLK 
            //to compensate for temperature and voltage variations.
            RXDLYEN[MASTER_LANE_ID] <= `DLY  1'b1;
            PHASE_ALIGNMENT_DONE    <= `DLY  1'b1;
           end

           default:
              rx_phalign_manual_state <= `DLY  INIT;

        endcase
      end 
    end   


endmodule

//------------------------------------------------------------------------------
//   ____  ____
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 3.5
//  \   \         Application : 7 Series FPGAs Transceivers Wizard 
//  /   /         Filename : gtwizard_0_init.v
// /___/   /\      
// \   \  /  \ 
//  \___\/\___\
//
//  Description : This module instantiates the modules required for
//                reset and initialisation of the Transceiver
//
// Module gtwizard_0_init
// Generated by Xilinx 7 Series FPGAs Transceivers Wizard
// 
// 
// (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES. 


`timescale 1ns / 1ps
`define DLY #1

//***********************************Entity Declaration************************
(* DowngradeIPIdentifiedWarnings="yes" *)
module gtwizard_0_init #
(
    parameter EXAMPLE_SIM_GTRESET_SPEEDUP            = "TRUE",     // Simulation setting for GT SecureIP model
    parameter EXAMPLE_SIMULATION                     =  0,         // Set to 1 for simulation
    parameter STABLE_CLOCK_PERIOD                    = 10,         //Period of the stable clock driving this state-machine, unit is [ns]
    parameter EXAMPLE_USE_CHIPSCOPE                  =  0          // Set to 1 to use Chipscope to drive resets

)
(
input           sysclk_in,
input           soft_reset_tx_in,
input           soft_reset_rx_in,
input           dont_reset_on_data_error_in,
output          gt0_tx_fsm_reset_done_out,
output          gt0_rx_fsm_reset_done_out,
input           gt0_data_valid_in,
output          gt1_tx_fsm_reset_done_out,
output          gt1_rx_fsm_reset_done_out,
input           gt1_data_valid_in,
output          gt2_tx_fsm_reset_done_out,
output          gt2_rx_fsm_reset_done_out,
input           gt2_data_valid_in,
output          gt3_tx_fsm_reset_done_out,
output          gt3_rx_fsm_reset_done_out,
input           gt3_data_valid_in,

    //_________________________________________________________________________
    //GT0  (X1Y4)
    //____________________________CHANNEL PORTS________________________________
    //------------------------ Channel - Clocking Ports ------------------------
    input           gt0_gtgrefclk_in,
    input           gt0_gtnorthrefclk0_in,
    input           gt0_gtnorthrefclk1_in,
    input           gt0_gtsouthrefclk0_in,
    input           gt0_gtsouthrefclk1_in,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt0_drpaddr_in,
    input           gt0_drpclk_in,
    input   [15:0]  gt0_drpdi_in,
    output  [15:0]  gt0_drpdo_out,
    input           gt0_drpen_in,
    output          gt0_drprdy_out,
    input           gt0_drpwe_in,
    //----------------------------- Clocking Ports -----------------------------
    input   [1:0]   gt0_txsysclksel_in,
    //------------------------- Digital Monitor Ports --------------------------
    output  [7:0]   gt0_dmonitorout_out,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   gt0_loopback_in,
    //--------------------------- PCI Express Ports ----------------------------
    input   [2:0]   gt0_rxrate_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt0_eyescanreset_in,
    input           gt0_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt0_eyescandataerror_out,
    input           gt0_eyescantrigger_in,
    //----------------------- Receive Ports - CDR Ports ------------------------
    input           gt0_rxcdrhold_in,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt0_rxusrclk_in,
    input           gt0_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [19:0]  gt0_rxdata_out,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           gt0_gtxrxp_in,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt0_gtxrxn_in,
    //----------------- Receive Ports - RX Buffer Bypass Ports -----------------
    input           gt0_rxbufreset_in,
    output  [2:0]   gt0_rxbufstatus_out,
    output  [4:0]   gt0_rxphmonitor_out,
    output  [4:0]   gt0_rxphslipmonitor_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    input           gt0_rxdfelpmreset_in,
    output  [6:0]   gt0_rxmonitorout_out,
    input   [1:0]   gt0_rxmonitorsel_in,
    //---------- Receive Ports - RX Fabric ClocK Output Control Ports ----------
    output          gt0_rxratedone_out,
    //------------- Receive Ports - RX Fabric Output Control Ports -------------
    output          gt0_rxoutclk_out,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt0_gtrxreset_in,
    input           gt0_rxpcsreset_in,
    input           gt0_rxpmareset_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt0_rxresetdone_out,
    //---------------------- TX Configurable Driver Ports ----------------------
    input   [4:0]   gt0_txpostcursor_in,
    input   [4:0]   gt0_txprecursor_in,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt0_gttxreset_in,
    input           gt0_txuserrdy_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt0_txusrclk_in,
    input           gt0_txusrclk2_in,
    //------------------- Transmit Ports - PCI Express Ports -------------------
    input   [2:0]   gt0_txrate_in,
    //-------------------- Transmit Ports - TX Buffer Ports --------------------
    output  [1:0]   gt0_txbufstatus_out,
    //------------- Transmit Ports - TX Configurable Driver Ports --------------
    input   [3:0]   gt0_txdiffctrl_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [19:0]  gt0_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt0_gtxtxn_out,
    output          gt0_gtxtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt0_txoutclk_out,
    output          gt0_txoutclkfabric_out,
    output          gt0_txoutclkpcs_out,
    output          gt0_txratedone_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    input           gt0_txpcsreset_in,
    input           gt0_txpmareset_in,
    output          gt0_txresetdone_out,

    //GT1  (X1Y5)
    //____________________________CHANNEL PORTS________________________________
    //------------------------ Channel - Clocking Ports ------------------------
    input           gt1_gtgrefclk_in,
    input           gt1_gtnorthrefclk0_in,
    input           gt1_gtnorthrefclk1_in,
    input           gt1_gtsouthrefclk0_in,
    input           gt1_gtsouthrefclk1_in,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt1_drpaddr_in,
    input           gt1_drpclk_in,
    input   [15:0]  gt1_drpdi_in,
    output  [15:0]  gt1_drpdo_out,
    input           gt1_drpen_in,
    output          gt1_drprdy_out,
    input           gt1_drpwe_in,
    //----------------------------- Clocking Ports -----------------------------
    input   [1:0]   gt1_txsysclksel_in,
    //------------------------- Digital Monitor Ports --------------------------
    output  [7:0]   gt1_dmonitorout_out,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   gt1_loopback_in,
    //--------------------------- PCI Express Ports ----------------------------
    input   [2:0]   gt1_rxrate_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt1_eyescanreset_in,
    input           gt1_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt1_eyescandataerror_out,
    input           gt1_eyescantrigger_in,
    //----------------------- Receive Ports - CDR Ports ------------------------
    input           gt1_rxcdrhold_in,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt1_rxusrclk_in,
    input           gt1_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [19:0]  gt1_rxdata_out,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           gt1_gtxrxp_in,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt1_gtxrxn_in,
    //----------------- Receive Ports - RX Buffer Bypass Ports -----------------
    input           gt1_rxbufreset_in,
    output  [2:0]   gt1_rxbufstatus_out,
    output  [4:0]   gt1_rxphmonitor_out,
    output  [4:0]   gt1_rxphslipmonitor_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    input           gt1_rxdfelpmreset_in,
    output  [6:0]   gt1_rxmonitorout_out,
    input   [1:0]   gt1_rxmonitorsel_in,
    //---------- Receive Ports - RX Fabric ClocK Output Control Ports ----------
    output          gt1_rxratedone_out,
    //------------- Receive Ports - RX Fabric Output Control Ports -------------
    output          gt1_rxoutclk_out,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt1_gtrxreset_in,
    input           gt1_rxpcsreset_in,
    input           gt1_rxpmareset_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt1_rxresetdone_out,
    //---------------------- TX Configurable Driver Ports ----------------------
    input   [4:0]   gt1_txpostcursor_in,
    input   [4:0]   gt1_txprecursor_in,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt1_gttxreset_in,
    input           gt1_txuserrdy_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt1_txusrclk_in,
    input           gt1_txusrclk2_in,
    //------------------- Transmit Ports - PCI Express Ports -------------------
    input   [2:0]   gt1_txrate_in,
    //-------------------- Transmit Ports - TX Buffer Ports --------------------
    output  [1:0]   gt1_txbufstatus_out,
    //------------- Transmit Ports - TX Configurable Driver Ports --------------
    input   [3:0]   gt1_txdiffctrl_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [19:0]  gt1_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt1_gtxtxn_out,
    output          gt1_gtxtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt1_txoutclk_out,
    output          gt1_txoutclkfabric_out,
    output          gt1_txoutclkpcs_out,
    output          gt1_txratedone_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    input           gt1_txpcsreset_in,
    input           gt1_txpmareset_in,
    output          gt1_txresetdone_out,

    //GT2  (X1Y6)
    //____________________________CHANNEL PORTS________________________________
    //------------------------ Channel - Clocking Ports ------------------------
    input           gt2_gtgrefclk_in,
    input           gt2_gtnorthrefclk0_in,
    input           gt2_gtnorthrefclk1_in,
    input           gt2_gtsouthrefclk0_in,
    input           gt2_gtsouthrefclk1_in,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt2_drpaddr_in,
    input           gt2_drpclk_in,
    input   [15:0]  gt2_drpdi_in,
    output  [15:0]  gt2_drpdo_out,
    input           gt2_drpen_in,
    output          gt2_drprdy_out,
    input           gt2_drpwe_in,
    //----------------------------- Clocking Ports -----------------------------
    input   [1:0]   gt2_txsysclksel_in,
    //------------------------- Digital Monitor Ports --------------------------
    output  [7:0]   gt2_dmonitorout_out,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   gt2_loopback_in,
    //--------------------------- PCI Express Ports ----------------------------
    input   [2:0]   gt2_rxrate_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt2_eyescanreset_in,
    input           gt2_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt2_eyescandataerror_out,
    input           gt2_eyescantrigger_in,
    //----------------------- Receive Ports - CDR Ports ------------------------
    input           gt2_rxcdrhold_in,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt2_rxusrclk_in,
    input           gt2_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [19:0]  gt2_rxdata_out,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           gt2_gtxrxp_in,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt2_gtxrxn_in,
    //----------------- Receive Ports - RX Buffer Bypass Ports -----------------
    input           gt2_rxbufreset_in,
    output  [2:0]   gt2_rxbufstatus_out,
    output  [4:0]   gt2_rxphmonitor_out,
    output  [4:0]   gt2_rxphslipmonitor_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    input           gt2_rxdfelpmreset_in,
    output  [6:0]   gt2_rxmonitorout_out,
    input   [1:0]   gt2_rxmonitorsel_in,
    //---------- Receive Ports - RX Fabric ClocK Output Control Ports ----------
    output          gt2_rxratedone_out,
    //------------- Receive Ports - RX Fabric Output Control Ports -------------
    output          gt2_rxoutclk_out,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt2_gtrxreset_in,
    input           gt2_rxpcsreset_in,
    input           gt2_rxpmareset_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt2_rxresetdone_out,
    //---------------------- TX Configurable Driver Ports ----------------------
    input   [4:0]   gt2_txpostcursor_in,
    input   [4:0]   gt2_txprecursor_in,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt2_gttxreset_in,
    input           gt2_txuserrdy_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt2_txusrclk_in,
    input           gt2_txusrclk2_in,
    //------------------- Transmit Ports - PCI Express Ports -------------------
    input   [2:0]   gt2_txrate_in,
    //-------------------- Transmit Ports - TX Buffer Ports --------------------
    output  [1:0]   gt2_txbufstatus_out,
    //------------- Transmit Ports - TX Configurable Driver Ports --------------
    input   [3:0]   gt2_txdiffctrl_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [19:0]  gt2_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt2_gtxtxn_out,
    output          gt2_gtxtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt2_txoutclk_out,
    output          gt2_txoutclkfabric_out,
    output          gt2_txoutclkpcs_out,
    output          gt2_txratedone_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    input           gt2_txpcsreset_in,
    input           gt2_txpmareset_in,
    output          gt2_txresetdone_out,

    //GT3  (X1Y7)
    //____________________________CHANNEL PORTS________________________________
    //------------------------ Channel - Clocking Ports ------------------------
    input           gt3_gtgrefclk_in,
    input           gt3_gtnorthrefclk0_in,
    input           gt3_gtnorthrefclk1_in,
    input           gt3_gtsouthrefclk0_in,
    input           gt3_gtsouthrefclk1_in,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   gt3_drpaddr_in,
    input           gt3_drpclk_in,
    input   [15:0]  gt3_drpdi_in,
    output  [15:0]  gt3_drpdo_out,
    input           gt3_drpen_in,
    output          gt3_drprdy_out,
    input           gt3_drpwe_in,
    //----------------------------- Clocking Ports -----------------------------
    input   [1:0]   gt3_txsysclksel_in,
    //------------------------- Digital Monitor Ports --------------------------
    output  [7:0]   gt3_dmonitorout_out,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   gt3_loopback_in,
    //--------------------------- PCI Express Ports ----------------------------
    input   [2:0]   gt3_rxrate_in,
    //------------------- RX Initialization and Reset Ports --------------------
    input           gt3_eyescanreset_in,
    input           gt3_rxuserrdy_in,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          gt3_eyescandataerror_out,
    input           gt3_eyescantrigger_in,
    //----------------------- Receive Ports - CDR Ports ------------------------
    input           gt3_rxcdrhold_in,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           gt3_rxusrclk_in,
    input           gt3_rxusrclk2_in,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [19:0]  gt3_rxdata_out,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           gt3_gtxrxp_in,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           gt3_gtxrxn_in,
    //----------------- Receive Ports - RX Buffer Bypass Ports -----------------
    input           gt3_rxbufreset_in,
    output  [2:0]   gt3_rxbufstatus_out,
    output  [4:0]   gt3_rxphmonitor_out,
    output  [4:0]   gt3_rxphslipmonitor_out,
    //------------------- Receive Ports - RX Equalizer Ports -------------------
    input           gt3_rxdfelpmreset_in,
    output  [6:0]   gt3_rxmonitorout_out,
    input   [1:0]   gt3_rxmonitorsel_in,
    //---------- Receive Ports - RX Fabric ClocK Output Control Ports ----------
    output          gt3_rxratedone_out,
    //------------- Receive Ports - RX Fabric Output Control Ports -------------
    output          gt3_rxoutclk_out,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           gt3_gtrxreset_in,
    input           gt3_rxpcsreset_in,
    input           gt3_rxpmareset_in,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          gt3_rxresetdone_out,
    //---------------------- TX Configurable Driver Ports ----------------------
    input   [4:0]   gt3_txpostcursor_in,
    input   [4:0]   gt3_txprecursor_in,
    //------------------- TX Initialization and Reset Ports --------------------
    input           gt3_gttxreset_in,
    input           gt3_txuserrdy_in,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           gt3_txusrclk_in,
    input           gt3_txusrclk2_in,
    //------------------- Transmit Ports - PCI Express Ports -------------------
    input   [2:0]   gt3_txrate_in,
    //-------------------- Transmit Ports - TX Buffer Ports --------------------
    output  [1:0]   gt3_txbufstatus_out,
    //------------- Transmit Ports - TX Configurable Driver Ports --------------
    input   [3:0]   gt3_txdiffctrl_in,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [19:0]  gt3_txdata_in,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          gt3_gtxtxn_out,
    output          gt3_gtxtxp_out,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          gt3_txoutclk_out,
    output          gt3_txoutclkfabric_out,
    output          gt3_txoutclkpcs_out,
    output          gt3_txratedone_out,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    input           gt3_txpcsreset_in,
    input           gt3_txpmareset_in,
    output          gt3_txresetdone_out,


    //____________________________COMMON PORTS________________________________
    input      gt0_qplllock_in,
    input      gt0_qpllrefclklost_in,
    output     gt0_qpllreset_out,
    input      gt0_qplloutclk_in,
    input      gt0_qplloutrefclk_in

);



//***********************************Parameter Declarations********************


    //Typical CDRLOCK Time is 50,000UI, as per DS183
    localparam RX_CDRLOCK_TIME      = (EXAMPLE_SIMULATION == 1) ? 1000 : 50000/2.97;
       
    integer   WAIT_TIME_CDRLOCK    = RX_CDRLOCK_TIME / STABLE_CLOCK_PERIOD;      

//-------------------------- GT Wrapper Wires ------------------------------
    wire           gt0_rxpmaresetdone_i;
    wire           gt0_txpmaresetdone_i;
    wire           gt0_txresetdone_i;
    wire           gt0_rxresetdone_i;
    wire           gt0_gttxreset_i;
    wire           gt0_gttxreset_t;
    wire           gt0_gtrxreset_i;
    wire           gt0_gtrxreset_t;
    wire           gt0_txpcsreset_i;
    wire           gt0_rxpcsreset_i;
    wire           gt0_txpmareset_i;
    wire           gt0_rxdfelpmreset_i;
    wire   [1:0]   gt0_txsysclksel_i;
    wire           gt0_txuserrdy_i;
    wire           gt0_txuserrdy_t;
    wire           gt0_rxuserrdy_i;
    wire           gt0_rxuserrdy_t;

    wire           gt0_rxdfeagchold_i;
    wire           gt0_rxdfelfhold_i;
    wire           gt0_rxlpmlfhold_i;
    wire           gt0_rxlpmhfhold_i;


    wire           gt1_rxpmaresetdone_i;
    wire           gt1_txpmaresetdone_i;
    wire           gt1_txresetdone_i;
    wire           gt1_rxresetdone_i;
    wire           gt1_gttxreset_i;
    wire           gt1_gttxreset_t;
    wire           gt1_gtrxreset_i;
    wire           gt1_gtrxreset_t;
    wire           gt1_txpcsreset_i;
    wire           gt1_rxpcsreset_i;
    wire           gt1_txpmareset_i;
    wire           gt1_rxdfelpmreset_i;
    wire   [1:0]   gt1_txsysclksel_i;
    wire           gt1_txuserrdy_i;
    wire           gt1_txuserrdy_t;
    wire           gt1_rxuserrdy_i;
    wire           gt1_rxuserrdy_t;

    wire           gt1_rxdfeagchold_i;
    wire           gt1_rxdfelfhold_i;
    wire           gt1_rxlpmlfhold_i;
    wire           gt1_rxlpmhfhold_i;


    wire           gt2_rxpmaresetdone_i;
    wire           gt2_txpmaresetdone_i;
    wire           gt2_txresetdone_i;
    wire           gt2_rxresetdone_i;
    wire           gt2_gttxreset_i;
    wire           gt2_gttxreset_t;
    wire           gt2_gtrxreset_i;
    wire           gt2_gtrxreset_t;
    wire           gt2_txpcsreset_i;
    wire           gt2_rxpcsreset_i;
    wire           gt2_txpmareset_i;
    wire           gt2_rxdfelpmreset_i;
    wire   [1:0]   gt2_txsysclksel_i;
    wire           gt2_txuserrdy_i;
    wire           gt2_txuserrdy_t;
    wire           gt2_rxuserrdy_i;
    wire           gt2_rxuserrdy_t;

    wire           gt2_rxdfeagchold_i;
    wire           gt2_rxdfelfhold_i;
    wire           gt2_rxlpmlfhold_i;
    wire           gt2_rxlpmhfhold_i;


    wire           gt3_rxpmaresetdone_i;
    wire           gt3_txpmaresetdone_i;
    wire           gt3_txresetdone_i;
    wire           gt3_rxresetdone_i;
    wire           gt3_gttxreset_i;
    wire           gt3_gttxreset_t;
    wire           gt3_gtrxreset_i;
    wire           gt3_gtrxreset_t;
    wire           gt3_txpcsreset_i;
    wire           gt3_rxpcsreset_i;
    wire           gt3_txpmareset_i;
    wire           gt3_rxdfelpmreset_i;
    wire   [1:0]   gt3_txsysclksel_i;
    wire           gt3_txuserrdy_i;
    wire           gt3_txuserrdy_t;
    wire           gt3_rxuserrdy_i;
    wire           gt3_rxuserrdy_t;

    wire           gt3_rxdfeagchold_i;
    wire           gt3_rxdfelfhold_i;
    wire           gt3_rxlpmlfhold_i;
    wire           gt3_rxlpmhfhold_i;



    wire           gt0_qpllreset_i;
    wire           gt0_qpllreset_t;
    wire           gt0_qpllrefclklost_i;
    wire           gt0_qplllock_i;


//------------------------------- Global Signals -----------------------------
    wire          tied_to_ground_i;
    wire          tied_to_vcc_i;
    wire           gt0_txphaligndone_i;
    wire           gt0_txdlysreset_i;
    wire           gt0_txdlysresetdone_i;
    wire           gt0_txphdlyreset_i;
    wire           gt0_txphalignen_i;
    wire           gt0_txdlyen_i;
    wire           gt0_txphalign_i;
    wire           gt0_txphinit_i;
    wire           gt0_txphinitdone_i;
    wire           gt0_run_tx_phalignment_i;
    wire           gt0_rst_tx_phalignment_i;
    wire           gt0_tx_phalignment_done_i;

    wire           gt0_txoutclk_i;
    wire           gt0_rxoutclk_i;
    wire           gt0_rxoutclk_i2;
    wire           gt0_txoutclk_i2;
    wire           gt0_recclk_stable_i;
    reg            gt0_rx_cdrlocked;
    integer  gt0_rx_cdrlock_counter= 0;
    wire           gt0_rxphaligndone_i;
    wire           gt0_rxdlysreset_i;
    wire           gt0_rxdlysresetdone_i;
    wire           gt0_rxphdlyreset_i;
    wire           gt0_rxphalignen_i;
    wire           gt0_rxdlyen_i;
    wire           gt0_rxphalign_i;
    wire           gt0_run_rx_phalignment_i;
    wire           gt0_rst_rx_phalignment_i;
    wire           gt0_rx_phalignment_done_i;
    wire           gt1_txphaligndone_i;
    wire           gt1_txdlysreset_i;
    wire           gt1_txdlysresetdone_i;
    wire           gt1_txphdlyreset_i;
    wire           gt1_txphalignen_i;
    wire           gt1_txdlyen_i;
    wire           gt1_txphalign_i;
    wire           gt1_txphinit_i;
    wire           gt1_txphinitdone_i;
    wire           gt1_run_tx_phalignment_i;
    wire           gt1_rst_tx_phalignment_i;
    wire           gt1_tx_phalignment_done_i;

    wire           gt1_txoutclk_i;
    wire           gt1_rxoutclk_i;
    wire           gt1_rxoutclk_i2;
    wire           gt1_txoutclk_i2;
    wire           gt1_recclk_stable_i;
    reg            gt1_rx_cdrlocked;
    integer  gt1_rx_cdrlock_counter= 0;
    wire           gt1_rxphaligndone_i;
    wire           gt1_rxdlysreset_i;
    wire           gt1_rxdlysresetdone_i;
    wire           gt1_rxphdlyreset_i;
    wire           gt1_rxphalignen_i;
    wire           gt1_rxdlyen_i;
    wire           gt1_rxphalign_i;
    wire           gt1_run_rx_phalignment_i;
    wire           gt1_rst_rx_phalignment_i;
    wire           gt1_rx_phalignment_done_i;
    wire           gt2_txphaligndone_i;
    wire           gt2_txdlysreset_i;
    wire           gt2_txdlysresetdone_i;
    wire           gt2_txphdlyreset_i;
    wire           gt2_txphalignen_i;
    wire           gt2_txdlyen_i;
    wire           gt2_txphalign_i;
    wire           gt2_txphinit_i;
    wire           gt2_txphinitdone_i;
    wire           gt2_run_tx_phalignment_i;
    wire           gt2_rst_tx_phalignment_i;
    wire           gt2_tx_phalignment_done_i;

    wire           gt2_txoutclk_i;
    wire           gt2_rxoutclk_i;
    wire           gt2_rxoutclk_i2;
    wire           gt2_txoutclk_i2;
    wire           gt2_recclk_stable_i;
    reg            gt2_rx_cdrlocked;
    integer  gt2_rx_cdrlock_counter= 0;
    wire           gt2_rxphaligndone_i;
    wire           gt2_rxdlysreset_i;
    wire           gt2_rxdlysresetdone_i;
    wire           gt2_rxphdlyreset_i;
    wire           gt2_rxphalignen_i;
    wire           gt2_rxdlyen_i;
    wire           gt2_rxphalign_i;
    wire           gt2_run_rx_phalignment_i;
    wire           gt2_rst_rx_phalignment_i;
    wire           gt2_rx_phalignment_done_i;
    wire           gt3_txphaligndone_i;
    wire           gt3_txdlysreset_i;
    wire           gt3_txdlysresetdone_i;
    wire           gt3_txphdlyreset_i;
    wire           gt3_txphalignen_i;
    wire           gt3_txdlyen_i;
    wire           gt3_txphalign_i;
    wire           gt3_txphinit_i;
    wire           gt3_txphinitdone_i;
    wire           gt3_run_tx_phalignment_i;
    wire           gt3_rst_tx_phalignment_i;
    wire           gt3_tx_phalignment_done_i;

    wire           gt3_txoutclk_i;
    wire           gt3_rxoutclk_i;
    wire           gt3_rxoutclk_i2;
    wire           gt3_txoutclk_i2;
    wire           gt3_recclk_stable_i;
    reg            gt3_rx_cdrlocked;
    integer  gt3_rx_cdrlock_counter= 0;
    wire           gt3_rxphaligndone_i;
    wire           gt3_rxdlysreset_i;
    wire           gt3_rxdlysresetdone_i;
    wire           gt3_rxphdlyreset_i;
    wire           gt3_rxphalignen_i;
    wire           gt3_rxdlyen_i;
    wire           gt3_rxphalign_i;
    wire           gt3_run_rx_phalignment_i;
    wire           gt3_rst_rx_phalignment_i;
    wire           gt3_rx_phalignment_done_i;



//    --------------------------- TX Buffer Bypass Signals --------------------
    wire   mstr0_txsyncallin_i;
    wire  [3 : 0]        U0_TXDLYEN;
    wire  [3 : 0]        U0_TXDLYSRESET;
    wire  [3 : 0]        U0_TXDLYSRESETDONE;
    wire  [3 : 0]        U0_TXPHINIT;
    wire  [3 : 0]        U0_TXPHINITDONE;
    wire  [3 : 0]        U0_TXPHALIGN;
    wire  [3 : 0]        U0_TXPHALIGNDONE ;
    wire                                 U0_run_tx_phalignment_i;
    wire                                 U0_rst_tx_phalignment_i;


//    --------------------------- RX Buffer Bypass Signals --------------------
    wire   rxmstr0_rxsyncallin_i;
    wire  [3 : 0]        U0_RXDLYEN;
    wire  [3 : 0]        U0_RXDLYSRESET;
    wire  [3 : 0]        U0_RXDLYSRESETDONE;
    wire  [3 : 0]        U0_RXPHALIGN;
    wire  [3 : 0]        U0_RXPHALIGNDONE ;
    wire                                 U0_run_rx_phalignment_i;
    wire                                 U0_rst_rx_phalignment_i;




reg              rx_cdrlocked;


 


//**************************** Main Body of Code *******************************
    //  Static signal Assigments
assign  tied_to_ground_i                     =  1'b0;
assign  tied_to_vcc_i                        =  1'b1;

//    ----------------------------- The GT Wrapper -----------------------------
    
    // Use the instantiation template in the example directory to add the GT wrapper to your design.
    // In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    // checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    // enabled, bonding should occur after alignment.


    gtwizard_0_multi_gt #
    (
        .WRAPPER_SIM_GTRESET_SPEEDUP    (EXAMPLE_SIM_GTRESET_SPEEDUP)
    )
    gtwizard_0_i
    (
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT0  (X1Y4)

        //------------------------ Channel - Clocking Ports ------------------------
        .gt0_gtgrefclk_in               (gt0_gtgrefclk_in), // input wire gt0_gtgrefclk_in
        .gt0_gtnorthrefclk0_in          (gt0_gtnorthrefclk0_in), // input wire gt0_gtnorthrefclk0_in
        .gt0_gtnorthrefclk1_in          (gt0_gtnorthrefclk1_in), // input wire gt0_gtnorthrefclk1_in
        .gt0_gtsouthrefclk0_in          (gt0_gtsouthrefclk0_in), // input wire gt0_gtsouthrefclk0_in
        .gt0_gtsouthrefclk1_in          (gt0_gtsouthrefclk1_in), // input wire gt0_gtsouthrefclk1_in
        //-------------------------- Channel - DRP Ports  --------------------------
        .gt0_drpaddr_in                 (gt0_drpaddr_in), // input wire [8:0] gt0_drpaddr_in
        .gt0_drpclk_in                  (gt0_drpclk_in), // input wire gt0_drpclk_in
        .gt0_drpdi_in                   (gt0_drpdi_in), // input wire [15:0] gt0_drpdi_in
        .gt0_drpdo_out                  (gt0_drpdo_out), // output wire [15:0] gt0_drpdo_out
        .gt0_drpen_in                   (gt0_drpen_in), // input wire gt0_drpen_in
        .gt0_drprdy_out                 (gt0_drprdy_out), // output wire gt0_drprdy_out
        .gt0_drpwe_in                   (gt0_drpwe_in), // input wire gt0_drpwe_in
        //----------------------------- Clocking Ports -----------------------------
        .gt0_txsysclksel_in             (gt0_txsysclksel_in), // input wire [1:0] gt0_txsysclksel_in
        //------------------------- Digital Monitor Ports --------------------------
        .gt0_dmonitorout_out            (gt0_dmonitorout_out), // output wire [7:0] gt0_dmonitorout_out
        //----------------------------- Loopback Ports -----------------------------
        .gt0_loopback_in                (gt0_loopback_in), // input wire [2:0] gt0_loopback_in
        //--------------------------- PCI Express Ports ----------------------------
        .gt0_rxrate_in                  (gt0_rxrate_in), // input wire [2:0] gt0_rxrate_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt0_eyescanreset_in            (gt0_eyescanreset_in), // input wire gt0_eyescanreset_in
        .gt0_rxuserrdy_in               (gt0_rxuserrdy_i), // input wire gt0_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt0_eyescandataerror_out       (gt0_eyescandataerror_out), // output wire gt0_eyescandataerror_out
        .gt0_eyescantrigger_in          (gt0_eyescantrigger_in), // input wire gt0_eyescantrigger_in
        //----------------------- Receive Ports - CDR Ports ------------------------
        .gt0_rxcdrhold_in               (gt0_rxcdrhold_in), // input wire gt0_rxcdrhold_in
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt0_rxusrclk_in                (gt0_rxusrclk_in), // input wire gt0_rxusrclk_in
        .gt0_rxusrclk2_in               (gt0_rxusrclk2_in), // input wire gt0_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt0_rxdata_out                 (gt0_rxdata_out), // output wire [19:0] gt0_rxdata_out
        //------------------------- Receive Ports - RX AFE -------------------------
        .gt0_gtxrxp_in                  (gt0_gtxrxp_in), // input wire gt0_gtxrxp_in
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt0_gtxrxn_in                  (gt0_gtxrxn_in), // input wire gt0_gtxrxn_in
        //----------------- Receive Ports - RX Buffer Bypass Ports -----------------
        .gt0_rxbufreset_in              (gt0_rxbufreset_in), // input wire gt0_rxbufreset_in
        .gt0_rxbufstatus_out            (gt0_rxbufstatus_out), // output wire [2:0] gt0_rxbufstatus_out
        .gt0_rxdlyen_in                 (gt0_rxdlyen_i), // input wire gt0_rxdlyen_i
        .gt0_rxdlysreset_in             (gt0_rxdlysreset_i), // input wire gt0_rxdlysreset_i
        .gt0_rxdlysresetdone_out        (gt0_rxdlysresetdone_i), // output wire gt0_rxdlysresetdone_i
        .gt0_rxphalign_in               (gt0_rxphalign_i), // input wire gt0_rxphalign_i
        .gt0_rxphaligndone_out          (gt0_rxphaligndone_i), // output wire gt0_rxphaligndone_i
        .gt0_rxphalignen_in             (gt0_rxphalignen_i), // input wire gt0_rxphalignen_i
        .gt0_rxphdlyreset_in            (gt0_rxphdlyreset_i), // input wire gt0_rxphdlyreset_i
        .gt0_rxphmonitor_out            (gt0_rxphmonitor_out), // output wire [4:0] gt0_rxphmonitor_out
        .gt0_rxphslipmonitor_out        (gt0_rxphslipmonitor_out), // output wire [4:0] gt0_rxphslipmonitor_out
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .gt0_rxlpmhfhold_in             (gt0_rxlpmhfhold_i), // input wire gt0_rxlpmhfhold_i
        .gt0_rxlpmlfhold_in             (gt0_rxlpmlfhold_i), // input wire gt0_rxlpmlfhold_i
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt0_rxdfelpmreset_in           (gt0_rxdfelpmreset_in), // input wire gt0_rxdfelpmreset_in
        .gt0_rxmonitorout_out           (gt0_rxmonitorout_out), // output wire [6:0] gt0_rxmonitorout_out
        .gt0_rxmonitorsel_in            (gt0_rxmonitorsel_in), // input wire [1:0] gt0_rxmonitorsel_in
        //---------- Receive Ports - RX Fabric ClocK Output Control Ports ----------
        .gt0_rxratedone_out             (gt0_rxratedone_out), // output wire gt0_rxratedone_out
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt0_rxoutclk_out               (gt0_rxoutclk_i), // output wire gt0_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt0_gtrxreset_in               (gt0_gtrxreset_i), // input wire gt0_gtrxreset_i
        .gt0_rxpcsreset_in              (gt0_rxpcsreset_in), // input wire gt0_rxpcsreset_in
        .gt0_rxpmareset_in              (gt0_rxpmareset_in), // input wire gt0_rxpmareset_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt0_rxresetdone_out            (gt0_rxresetdone_i), // output wire gt0_rxresetdone_i
        //---------------------- TX Configurable Driver Ports ----------------------
        .gt0_txpostcursor_in            (gt0_txpostcursor_in), // input wire [4:0] gt0_txpostcursor_in
        .gt0_txprecursor_in             (gt0_txprecursor_in), // input wire [4:0] gt0_txprecursor_in
        //------------------- TX Initialization and Reset Ports --------------------
        .gt0_gttxreset_in               (gt0_gttxreset_i), // input wire gt0_gttxreset_i
        .gt0_txuserrdy_in               (gt0_txuserrdy_i), // input wire gt0_txuserrdy_i
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt0_txusrclk_in                (gt0_txusrclk_in), // input wire gt0_txusrclk_in
        .gt0_txusrclk2_in               (gt0_txusrclk2_in), // input wire gt0_txusrclk2_in
        //------------------- Transmit Ports - PCI Express Ports -------------------
        .gt0_txrate_in                  (gt0_txrate_in), // input wire [2:0] gt0_txrate_in
        //---------------- Transmit Ports - TX Buffer Bypass Ports -----------------
        .gt0_txdlyen_in                 (gt0_txdlyen_i), // input wire gt0_txdlyen_i
        .gt0_txdlysreset_in             (gt0_txdlysreset_i), // input wire gt0_txdlysreset_i
        .gt0_txdlysresetdone_out        (gt0_txdlysresetdone_i), // output wire gt0_txdlysresetdone_i
        .gt0_txphalign_in               (gt0_txphalign_i), // input wire gt0_txphalign_i
        .gt0_txphaligndone_out          (gt0_txphaligndone_i), // output wire gt0_txphaligndone_i
        .gt0_txphalignen_in             (gt0_txphalignen_i), // input wire gt0_txphalignen_i
        .gt0_txphdlyreset_in            (gt0_txphdlyreset_i), // input wire gt0_txphdlyreset_i
        .gt0_txphinit_in                (gt0_txphinit_i), // input wire gt0_txphinit_i
        .gt0_txphinitdone_out           (gt0_txphinitdone_i), // output wire gt0_txphinitdone_i
        //-------------------- Transmit Ports - TX Buffer Ports --------------------
        .gt0_txbufstatus_out            (gt0_txbufstatus_out), // output wire [1:0] gt0_txbufstatus_out
        //------------- Transmit Ports - TX Configurable Driver Ports --------------
        .gt0_txdiffctrl_in              (gt0_txdiffctrl_in), // input wire [3:0] gt0_txdiffctrl_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt0_txdata_in                  (gt0_txdata_in), // input wire [19:0] gt0_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt0_gtxtxn_out                 (gt0_gtxtxn_out), // output wire gt0_gtxtxn_out
        .gt0_gtxtxp_out                 (gt0_gtxtxp_out), // output wire gt0_gtxtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt0_txoutclk_out               (gt0_txoutclk_i), // output wire gt0_txoutclk_i
        .gt0_txoutclkfabric_out         (gt0_txoutclkfabric_out), // output wire gt0_txoutclkfabric_out
        .gt0_txoutclkpcs_out            (gt0_txoutclkpcs_out), // output wire gt0_txoutclkpcs_out
        .gt0_txratedone_out             (gt0_txratedone_out), // output wire gt0_txratedone_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt0_txpcsreset_in              (gt0_txpcsreset_in), // input wire gt0_txpcsreset_in
        .gt0_txpmareset_in              (gt0_txpmareset_in), // input wire gt0_txpmareset_in
        .gt0_txresetdone_out            (gt0_txresetdone_i), // output wire gt0_txresetdone_i


 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT1  (X1Y5)

        //------------------------ Channel - Clocking Ports ------------------------
        .gt1_gtgrefclk_in               (gt1_gtgrefclk_in), // input wire gt1_gtgrefclk_in
        .gt1_gtnorthrefclk0_in          (gt1_gtnorthrefclk0_in), // input wire gt1_gtnorthrefclk0_in
        .gt1_gtnorthrefclk1_in          (gt1_gtnorthrefclk1_in), // input wire gt1_gtnorthrefclk1_in
        .gt1_gtsouthrefclk0_in          (gt1_gtsouthrefclk0_in), // input wire gt1_gtsouthrefclk0_in
        .gt1_gtsouthrefclk1_in          (gt1_gtsouthrefclk1_in), // input wire gt1_gtsouthrefclk1_in
        //-------------------------- Channel - DRP Ports  --------------------------
        .gt1_drpaddr_in                 (gt1_drpaddr_in), // input wire [8:0] gt1_drpaddr_in
        .gt1_drpclk_in                  (gt1_drpclk_in), // input wire gt1_drpclk_in
        .gt1_drpdi_in                   (gt1_drpdi_in), // input wire [15:0] gt1_drpdi_in
        .gt1_drpdo_out                  (gt1_drpdo_out), // output wire [15:0] gt1_drpdo_out
        .gt1_drpen_in                   (gt1_drpen_in), // input wire gt1_drpen_in
        .gt1_drprdy_out                 (gt1_drprdy_out), // output wire gt1_drprdy_out
        .gt1_drpwe_in                   (gt1_drpwe_in), // input wire gt1_drpwe_in
        //----------------------------- Clocking Ports -----------------------------
        .gt1_txsysclksel_in             (gt1_txsysclksel_in), // input wire [1:0] gt1_txsysclksel_in
        //------------------------- Digital Monitor Ports --------------------------
        .gt1_dmonitorout_out            (gt1_dmonitorout_out), // output wire [7:0] gt1_dmonitorout_out
        //----------------------------- Loopback Ports -----------------------------
        .gt1_loopback_in                (gt1_loopback_in), // input wire [2:0] gt1_loopback_in
        //--------------------------- PCI Express Ports ----------------------------
        .gt1_rxrate_in                  (gt1_rxrate_in), // input wire [2:0] gt1_rxrate_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt1_eyescanreset_in            (gt1_eyescanreset_in), // input wire gt1_eyescanreset_in
        .gt1_rxuserrdy_in               (gt1_rxuserrdy_i), // input wire gt1_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt1_eyescandataerror_out       (gt1_eyescandataerror_out), // output wire gt1_eyescandataerror_out
        .gt1_eyescantrigger_in          (gt1_eyescantrigger_in), // input wire gt1_eyescantrigger_in
        //----------------------- Receive Ports - CDR Ports ------------------------
        .gt1_rxcdrhold_in               (gt1_rxcdrhold_in), // input wire gt1_rxcdrhold_in
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt1_rxusrclk_in                (gt1_rxusrclk_in), // input wire gt1_rxusrclk_in
        .gt1_rxusrclk2_in               (gt1_rxusrclk2_in), // input wire gt1_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt1_rxdata_out                 (gt1_rxdata_out), // output wire [19:0] gt1_rxdata_out
        //------------------------- Receive Ports - RX AFE -------------------------
        .gt1_gtxrxp_in                  (gt1_gtxrxp_in), // input wire gt1_gtxrxp_in
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt1_gtxrxn_in                  (gt1_gtxrxn_in), // input wire gt1_gtxrxn_in
        //----------------- Receive Ports - RX Buffer Bypass Ports -----------------
        .gt1_rxbufreset_in              (gt1_rxbufreset_in), // input wire gt1_rxbufreset_in
        .gt1_rxbufstatus_out            (gt1_rxbufstatus_out), // output wire [2:0] gt1_rxbufstatus_out
        .gt1_rxdlyen_in                 (gt1_rxdlyen_i), // input wire gt1_rxdlyen_i
        .gt1_rxdlysreset_in             (gt1_rxdlysreset_i), // input wire gt1_rxdlysreset_i
        .gt1_rxdlysresetdone_out        (gt1_rxdlysresetdone_i), // output wire gt1_rxdlysresetdone_i
        .gt1_rxphalign_in               (gt1_rxphalign_i), // input wire gt1_rxphalign_i
        .gt1_rxphaligndone_out          (gt1_rxphaligndone_i), // output wire gt1_rxphaligndone_i
        .gt1_rxphalignen_in             (gt1_rxphalignen_i), // input wire gt1_rxphalignen_i
        .gt1_rxphdlyreset_in            (gt1_rxphdlyreset_i), // input wire gt1_rxphdlyreset_i
        .gt1_rxphmonitor_out            (gt1_rxphmonitor_out), // output wire [4:0] gt1_rxphmonitor_out
        .gt1_rxphslipmonitor_out        (gt1_rxphslipmonitor_out), // output wire [4:0] gt1_rxphslipmonitor_out
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .gt1_rxlpmhfhold_in             (gt1_rxlpmhfhold_i), // input wire gt1_rxlpmhfhold_i
        .gt1_rxlpmlfhold_in             (gt1_rxlpmlfhold_i), // input wire gt1_rxlpmlfhold_i
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt1_rxdfelpmreset_in           (gt1_rxdfelpmreset_in), // input wire gt1_rxdfelpmreset_in
        .gt1_rxmonitorout_out           (gt1_rxmonitorout_out), // output wire [6:0] gt1_rxmonitorout_out
        .gt1_rxmonitorsel_in            (gt1_rxmonitorsel_in), // input wire [1:0] gt1_rxmonitorsel_in
        //---------- Receive Ports - RX Fabric ClocK Output Control Ports ----------
        .gt1_rxratedone_out             (gt1_rxratedone_out), // output wire gt1_rxratedone_out
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt1_rxoutclk_out               (gt1_rxoutclk_i), // output wire gt1_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt1_gtrxreset_in               (gt1_gtrxreset_i), // input wire gt1_gtrxreset_i
        .gt1_rxpcsreset_in              (gt1_rxpcsreset_in), // input wire gt1_rxpcsreset_in
        .gt1_rxpmareset_in              (gt1_rxpmareset_in), // input wire gt1_rxpmareset_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt1_rxresetdone_out            (gt1_rxresetdone_i), // output wire gt1_rxresetdone_i
        //---------------------- TX Configurable Driver Ports ----------------------
        .gt1_txpostcursor_in            (gt1_txpostcursor_in), // input wire [4:0] gt1_txpostcursor_in
        .gt1_txprecursor_in             (gt1_txprecursor_in), // input wire [4:0] gt1_txprecursor_in
        //------------------- TX Initialization and Reset Ports --------------------
        .gt1_gttxreset_in               (gt1_gttxreset_i), // input wire gt1_gttxreset_i
        .gt1_txuserrdy_in               (gt1_txuserrdy_i), // input wire gt1_txuserrdy_i
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt1_txusrclk_in                (gt1_txusrclk_in), // input wire gt1_txusrclk_in
        .gt1_txusrclk2_in               (gt1_txusrclk2_in), // input wire gt1_txusrclk2_in
        //------------------- Transmit Ports - PCI Express Ports -------------------
        .gt1_txrate_in                  (gt1_txrate_in), // input wire [2:0] gt1_txrate_in
        //---------------- Transmit Ports - TX Buffer Bypass Ports -----------------
        .gt1_txdlyen_in                 (gt1_txdlyen_i), // input wire gt1_txdlyen_i
        .gt1_txdlysreset_in             (gt1_txdlysreset_i), // input wire gt1_txdlysreset_i
        .gt1_txdlysresetdone_out        (gt1_txdlysresetdone_i), // output wire gt1_txdlysresetdone_i
        .gt1_txphalign_in               (gt1_txphalign_i), // input wire gt1_txphalign_i
        .gt1_txphaligndone_out          (gt1_txphaligndone_i), // output wire gt1_txphaligndone_i
        .gt1_txphalignen_in             (gt1_txphalignen_i), // input wire gt1_txphalignen_i
        .gt1_txphdlyreset_in            (gt1_txphdlyreset_i), // input wire gt1_txphdlyreset_i
        .gt1_txphinit_in                (gt1_txphinit_i), // input wire gt1_txphinit_i
        .gt1_txphinitdone_out           (gt1_txphinitdone_i), // output wire gt1_txphinitdone_i
        //-------------------- Transmit Ports - TX Buffer Ports --------------------
        .gt1_txbufstatus_out            (gt1_txbufstatus_out), // output wire [1:0] gt1_txbufstatus_out
        //------------- Transmit Ports - TX Configurable Driver Ports --------------
        .gt1_txdiffctrl_in              (gt1_txdiffctrl_in), // input wire [3:0] gt1_txdiffctrl_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt1_txdata_in                  (gt1_txdata_in), // input wire [19:0] gt1_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt1_gtxtxn_out                 (gt1_gtxtxn_out), // output wire gt1_gtxtxn_out
        .gt1_gtxtxp_out                 (gt1_gtxtxp_out), // output wire gt1_gtxtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt1_txoutclk_out               (gt1_txoutclk_i), // output wire gt1_txoutclk_i
        .gt1_txoutclkfabric_out         (gt1_txoutclkfabric_out), // output wire gt1_txoutclkfabric_out
        .gt1_txoutclkpcs_out            (gt1_txoutclkpcs_out), // output wire gt1_txoutclkpcs_out
        .gt1_txratedone_out             (gt1_txratedone_out), // output wire gt1_txratedone_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt1_txpcsreset_in              (gt1_txpcsreset_in), // input wire gt1_txpcsreset_in
        .gt1_txpmareset_in              (gt1_txpmareset_in), // input wire gt1_txpmareset_in
        .gt1_txresetdone_out            (gt1_txresetdone_i), // output wire gt1_txresetdone_i


 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT2  (X1Y6)

        //------------------------ Channel - Clocking Ports ------------------------
        .gt2_gtgrefclk_in               (gt2_gtgrefclk_in), // input wire gt2_gtgrefclk_in
        .gt2_gtnorthrefclk0_in          (gt2_gtnorthrefclk0_in), // input wire gt2_gtnorthrefclk0_in
        .gt2_gtnorthrefclk1_in          (gt2_gtnorthrefclk1_in), // input wire gt2_gtnorthrefclk1_in
        .gt2_gtsouthrefclk0_in          (gt2_gtsouthrefclk0_in), // input wire gt2_gtsouthrefclk0_in
        .gt2_gtsouthrefclk1_in          (gt2_gtsouthrefclk1_in), // input wire gt2_gtsouthrefclk1_in
        //-------------------------- Channel - DRP Ports  --------------------------
        .gt2_drpaddr_in                 (gt2_drpaddr_in), // input wire [8:0] gt2_drpaddr_in
        .gt2_drpclk_in                  (gt2_drpclk_in), // input wire gt2_drpclk_in
        .gt2_drpdi_in                   (gt2_drpdi_in), // input wire [15:0] gt2_drpdi_in
        .gt2_drpdo_out                  (gt2_drpdo_out), // output wire [15:0] gt2_drpdo_out
        .gt2_drpen_in                   (gt2_drpen_in), // input wire gt2_drpen_in
        .gt2_drprdy_out                 (gt2_drprdy_out), // output wire gt2_drprdy_out
        .gt2_drpwe_in                   (gt2_drpwe_in), // input wire gt2_drpwe_in
        //----------------------------- Clocking Ports -----------------------------
        .gt2_txsysclksel_in             (gt2_txsysclksel_in), // input wire [1:0] gt2_txsysclksel_in
        //------------------------- Digital Monitor Ports --------------------------
        .gt2_dmonitorout_out            (gt2_dmonitorout_out), // output wire [7:0] gt2_dmonitorout_out
        //----------------------------- Loopback Ports -----------------------------
        .gt2_loopback_in                (gt2_loopback_in), // input wire [2:0] gt2_loopback_in
        //--------------------------- PCI Express Ports ----------------------------
        .gt2_rxrate_in                  (gt2_rxrate_in), // input wire [2:0] gt2_rxrate_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt2_eyescanreset_in            (gt2_eyescanreset_in), // input wire gt2_eyescanreset_in
        .gt2_rxuserrdy_in               (gt2_rxuserrdy_i), // input wire gt2_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt2_eyescandataerror_out       (gt2_eyescandataerror_out), // output wire gt2_eyescandataerror_out
        .gt2_eyescantrigger_in          (gt2_eyescantrigger_in), // input wire gt2_eyescantrigger_in
        //----------------------- Receive Ports - CDR Ports ------------------------
        .gt2_rxcdrhold_in               (gt2_rxcdrhold_in), // input wire gt2_rxcdrhold_in
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt2_rxusrclk_in                (gt2_rxusrclk_in), // input wire gt2_rxusrclk_in
        .gt2_rxusrclk2_in               (gt2_rxusrclk2_in), // input wire gt2_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt2_rxdata_out                 (gt2_rxdata_out), // output wire [19:0] gt2_rxdata_out
        //------------------------- Receive Ports - RX AFE -------------------------
        .gt2_gtxrxp_in                  (gt2_gtxrxp_in), // input wire gt2_gtxrxp_in
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt2_gtxrxn_in                  (gt2_gtxrxn_in), // input wire gt2_gtxrxn_in
        //----------------- Receive Ports - RX Buffer Bypass Ports -----------------
        .gt2_rxbufreset_in              (gt2_rxbufreset_in), // input wire gt2_rxbufreset_in
        .gt2_rxbufstatus_out            (gt2_rxbufstatus_out), // output wire [2:0] gt2_rxbufstatus_out
        .gt2_rxdlyen_in                 (gt2_rxdlyen_i), // input wire gt2_rxdlyen_i
        .gt2_rxdlysreset_in             (gt2_rxdlysreset_i), // input wire gt2_rxdlysreset_i
        .gt2_rxdlysresetdone_out        (gt2_rxdlysresetdone_i), // output wire gt2_rxdlysresetdone_i
        .gt2_rxphalign_in               (gt2_rxphalign_i), // input wire gt2_rxphalign_i
        .gt2_rxphaligndone_out          (gt2_rxphaligndone_i), // output wire gt2_rxphaligndone_i
        .gt2_rxphalignen_in             (gt2_rxphalignen_i), // input wire gt2_rxphalignen_i
        .gt2_rxphdlyreset_in            (gt2_rxphdlyreset_i), // input wire gt2_rxphdlyreset_i
        .gt2_rxphmonitor_out            (gt2_rxphmonitor_out), // output wire [4:0] gt2_rxphmonitor_out
        .gt2_rxphslipmonitor_out        (gt2_rxphslipmonitor_out), // output wire [4:0] gt2_rxphslipmonitor_out
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .gt2_rxlpmhfhold_in             (gt2_rxlpmhfhold_i), // input wire gt2_rxlpmhfhold_i
        .gt2_rxlpmlfhold_in             (gt2_rxlpmlfhold_i), // input wire gt2_rxlpmlfhold_i
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt2_rxdfelpmreset_in           (gt2_rxdfelpmreset_in), // input wire gt2_rxdfelpmreset_in
        .gt2_rxmonitorout_out           (gt2_rxmonitorout_out), // output wire [6:0] gt2_rxmonitorout_out
        .gt2_rxmonitorsel_in            (gt2_rxmonitorsel_in), // input wire [1:0] gt2_rxmonitorsel_in
        //---------- Receive Ports - RX Fabric ClocK Output Control Ports ----------
        .gt2_rxratedone_out             (gt2_rxratedone_out), // output wire gt2_rxratedone_out
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt2_rxoutclk_out               (gt2_rxoutclk_i), // output wire gt2_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt2_gtrxreset_in               (gt2_gtrxreset_i), // input wire gt2_gtrxreset_i
        .gt2_rxpcsreset_in              (gt2_rxpcsreset_in), // input wire gt2_rxpcsreset_in
        .gt2_rxpmareset_in              (gt2_rxpmareset_in), // input wire gt2_rxpmareset_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt2_rxresetdone_out            (gt2_rxresetdone_i), // output wire gt2_rxresetdone_i
        //---------------------- TX Configurable Driver Ports ----------------------
        .gt2_txpostcursor_in            (gt2_txpostcursor_in), // input wire [4:0] gt2_txpostcursor_in
        .gt2_txprecursor_in             (gt2_txprecursor_in), // input wire [4:0] gt2_txprecursor_in
        //------------------- TX Initialization and Reset Ports --------------------
        .gt2_gttxreset_in               (gt2_gttxreset_i), // input wire gt2_gttxreset_i
        .gt2_txuserrdy_in               (gt2_txuserrdy_i), // input wire gt2_txuserrdy_i
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt2_txusrclk_in                (gt2_txusrclk_in), // input wire gt2_txusrclk_in
        .gt2_txusrclk2_in               (gt2_txusrclk2_in), // input wire gt2_txusrclk2_in
        //------------------- Transmit Ports - PCI Express Ports -------------------
        .gt2_txrate_in                  (gt2_txrate_in), // input wire [2:0] gt2_txrate_in
        //---------------- Transmit Ports - TX Buffer Bypass Ports -----------------
        .gt2_txdlyen_in                 (gt2_txdlyen_i), // input wire gt2_txdlyen_i
        .gt2_txdlysreset_in             (gt2_txdlysreset_i), // input wire gt2_txdlysreset_i
        .gt2_txdlysresetdone_out        (gt2_txdlysresetdone_i), // output wire gt2_txdlysresetdone_i
        .gt2_txphalign_in               (gt2_txphalign_i), // input wire gt2_txphalign_i
        .gt2_txphaligndone_out          (gt2_txphaligndone_i), // output wire gt2_txphaligndone_i
        .gt2_txphalignen_in             (gt2_txphalignen_i), // input wire gt2_txphalignen_i
        .gt2_txphdlyreset_in            (gt2_txphdlyreset_i), // input wire gt2_txphdlyreset_i
        .gt2_txphinit_in                (gt2_txphinit_i), // input wire gt2_txphinit_i
        .gt2_txphinitdone_out           (gt2_txphinitdone_i), // output wire gt2_txphinitdone_i
        //-------------------- Transmit Ports - TX Buffer Ports --------------------
        .gt2_txbufstatus_out            (gt2_txbufstatus_out), // output wire [1:0] gt2_txbufstatus_out
        //------------- Transmit Ports - TX Configurable Driver Ports --------------
        .gt2_txdiffctrl_in              (gt2_txdiffctrl_in), // input wire [3:0] gt2_txdiffctrl_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt2_txdata_in                  (gt2_txdata_in), // input wire [19:0] gt2_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt2_gtxtxn_out                 (gt2_gtxtxn_out), // output wire gt2_gtxtxn_out
        .gt2_gtxtxp_out                 (gt2_gtxtxp_out), // output wire gt2_gtxtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt2_txoutclk_out               (gt2_txoutclk_i), // output wire gt2_txoutclk_i
        .gt2_txoutclkfabric_out         (gt2_txoutclkfabric_out), // output wire gt2_txoutclkfabric_out
        .gt2_txoutclkpcs_out            (gt2_txoutclkpcs_out), // output wire gt2_txoutclkpcs_out
        .gt2_txratedone_out             (gt2_txratedone_out), // output wire gt2_txratedone_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt2_txpcsreset_in              (gt2_txpcsreset_in), // input wire gt2_txpcsreset_in
        .gt2_txpmareset_in              (gt2_txpmareset_in), // input wire gt2_txpmareset_in
        .gt2_txresetdone_out            (gt2_txresetdone_i), // output wire gt2_txresetdone_i


 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT3  (X1Y7)

        //------------------------ Channel - Clocking Ports ------------------------
        .gt3_gtgrefclk_in               (gt3_gtgrefclk_in), // input wire gt3_gtgrefclk_in
        .gt3_gtnorthrefclk0_in          (gt3_gtnorthrefclk0_in), // input wire gt3_gtnorthrefclk0_in
        .gt3_gtnorthrefclk1_in          (gt3_gtnorthrefclk1_in), // input wire gt3_gtnorthrefclk1_in
        .gt3_gtsouthrefclk0_in          (gt3_gtsouthrefclk0_in), // input wire gt3_gtsouthrefclk0_in
        .gt3_gtsouthrefclk1_in          (gt3_gtsouthrefclk1_in), // input wire gt3_gtsouthrefclk1_in
        //-------------------------- Channel - DRP Ports  --------------------------
        .gt3_drpaddr_in                 (gt3_drpaddr_in), // input wire [8:0] gt3_drpaddr_in
        .gt3_drpclk_in                  (gt3_drpclk_in), // input wire gt3_drpclk_in
        .gt3_drpdi_in                   (gt3_drpdi_in), // input wire [15:0] gt3_drpdi_in
        .gt3_drpdo_out                  (gt3_drpdo_out), // output wire [15:0] gt3_drpdo_out
        .gt3_drpen_in                   (gt3_drpen_in), // input wire gt3_drpen_in
        .gt3_drprdy_out                 (gt3_drprdy_out), // output wire gt3_drprdy_out
        .gt3_drpwe_in                   (gt3_drpwe_in), // input wire gt3_drpwe_in
        //----------------------------- Clocking Ports -----------------------------
        .gt3_txsysclksel_in             (gt3_txsysclksel_in), // input wire [1:0] gt3_txsysclksel_in
        //------------------------- Digital Monitor Ports --------------------------
        .gt3_dmonitorout_out            (gt3_dmonitorout_out), // output wire [7:0] gt3_dmonitorout_out
        //----------------------------- Loopback Ports -----------------------------
        .gt3_loopback_in                (gt3_loopback_in), // input wire [2:0] gt3_loopback_in
        //--------------------------- PCI Express Ports ----------------------------
        .gt3_rxrate_in                  (gt3_rxrate_in), // input wire [2:0] gt3_rxrate_in
        //------------------- RX Initialization and Reset Ports --------------------
        .gt3_eyescanreset_in            (gt3_eyescanreset_in), // input wire gt3_eyescanreset_in
        .gt3_rxuserrdy_in               (gt3_rxuserrdy_i), // input wire gt3_rxuserrdy_i
        //------------------------ RX Margin Analysis Ports ------------------------
        .gt3_eyescandataerror_out       (gt3_eyescandataerror_out), // output wire gt3_eyescandataerror_out
        .gt3_eyescantrigger_in          (gt3_eyescantrigger_in), // input wire gt3_eyescantrigger_in
        //----------------------- Receive Ports - CDR Ports ------------------------
        .gt3_rxcdrhold_in               (gt3_rxcdrhold_in), // input wire gt3_rxcdrhold_in
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .gt3_rxusrclk_in                (gt3_rxusrclk_in), // input wire gt3_rxusrclk_in
        .gt3_rxusrclk2_in               (gt3_rxusrclk2_in), // input wire gt3_rxusrclk2_in
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .gt3_rxdata_out                 (gt3_rxdata_out), // output wire [19:0] gt3_rxdata_out
        //------------------------- Receive Ports - RX AFE -------------------------
        .gt3_gtxrxp_in                  (gt3_gtxrxp_in), // input wire gt3_gtxrxp_in
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .gt3_gtxrxn_in                  (gt3_gtxrxn_in), // input wire gt3_gtxrxn_in
        //----------------- Receive Ports - RX Buffer Bypass Ports -----------------
        .gt3_rxbufreset_in              (gt3_rxbufreset_in), // input wire gt3_rxbufreset_in
        .gt3_rxbufstatus_out            (gt3_rxbufstatus_out), // output wire [2:0] gt3_rxbufstatus_out
        .gt3_rxdlyen_in                 (gt3_rxdlyen_i), // input wire gt3_rxdlyen_i
        .gt3_rxdlysreset_in             (gt3_rxdlysreset_i), // input wire gt3_rxdlysreset_i
        .gt3_rxdlysresetdone_out        (gt3_rxdlysresetdone_i), // output wire gt3_rxdlysresetdone_i
        .gt3_rxphalign_in               (gt3_rxphalign_i), // input wire gt3_rxphalign_i
        .gt3_rxphaligndone_out          (gt3_rxphaligndone_i), // output wire gt3_rxphaligndone_i
        .gt3_rxphalignen_in             (gt3_rxphalignen_i), // input wire gt3_rxphalignen_i
        .gt3_rxphdlyreset_in            (gt3_rxphdlyreset_i), // input wire gt3_rxphdlyreset_i
        .gt3_rxphmonitor_out            (gt3_rxphmonitor_out), // output wire [4:0] gt3_rxphmonitor_out
        .gt3_rxphslipmonitor_out        (gt3_rxphslipmonitor_out), // output wire [4:0] gt3_rxphslipmonitor_out
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .gt3_rxlpmhfhold_in             (gt3_rxlpmhfhold_i), // input wire gt3_rxlpmhfhold_i
        .gt3_rxlpmlfhold_in             (gt3_rxlpmlfhold_i), // input wire gt3_rxlpmlfhold_i
        //------------------- Receive Ports - RX Equalizer Ports -------------------
        .gt3_rxdfelpmreset_in           (gt3_rxdfelpmreset_in), // input wire gt3_rxdfelpmreset_in
        .gt3_rxmonitorout_out           (gt3_rxmonitorout_out), // output wire [6:0] gt3_rxmonitorout_out
        .gt3_rxmonitorsel_in            (gt3_rxmonitorsel_in), // input wire [1:0] gt3_rxmonitorsel_in
        //---------- Receive Ports - RX Fabric ClocK Output Control Ports ----------
        .gt3_rxratedone_out             (gt3_rxratedone_out), // output wire gt3_rxratedone_out
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .gt3_rxoutclk_out               (gt3_rxoutclk_i), // output wire gt3_rxoutclk_i
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .gt3_gtrxreset_in               (gt3_gtrxreset_i), // input wire gt3_gtrxreset_i
        .gt3_rxpcsreset_in              (gt3_rxpcsreset_in), // input wire gt3_rxpcsreset_in
        .gt3_rxpmareset_in              (gt3_rxpmareset_in), // input wire gt3_rxpmareset_in
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .gt3_rxresetdone_out            (gt3_rxresetdone_i), // output wire gt3_rxresetdone_i
        //---------------------- TX Configurable Driver Ports ----------------------
        .gt3_txpostcursor_in            (gt3_txpostcursor_in), // input wire [4:0] gt3_txpostcursor_in
        .gt3_txprecursor_in             (gt3_txprecursor_in), // input wire [4:0] gt3_txprecursor_in
        //------------------- TX Initialization and Reset Ports --------------------
        .gt3_gttxreset_in               (gt3_gttxreset_i), // input wire gt3_gttxreset_i
        .gt3_txuserrdy_in               (gt3_txuserrdy_i), // input wire gt3_txuserrdy_i
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .gt3_txusrclk_in                (gt3_txusrclk_in), // input wire gt3_txusrclk_in
        .gt3_txusrclk2_in               (gt3_txusrclk2_in), // input wire gt3_txusrclk2_in
        //------------------- Transmit Ports - PCI Express Ports -------------------
        .gt3_txrate_in                  (gt3_txrate_in), // input wire [2:0] gt3_txrate_in
        //---------------- Transmit Ports - TX Buffer Bypass Ports -----------------
        .gt3_txdlyen_in                 (gt3_txdlyen_i), // input wire gt3_txdlyen_i
        .gt3_txdlysreset_in             (gt3_txdlysreset_i), // input wire gt3_txdlysreset_i
        .gt3_txdlysresetdone_out        (gt3_txdlysresetdone_i), // output wire gt3_txdlysresetdone_i
        .gt3_txphalign_in               (gt3_txphalign_i), // input wire gt3_txphalign_i
        .gt3_txphaligndone_out          (gt3_txphaligndone_i), // output wire gt3_txphaligndone_i
        .gt3_txphalignen_in             (gt3_txphalignen_i), // input wire gt3_txphalignen_i
        .gt3_txphdlyreset_in            (gt3_txphdlyreset_i), // input wire gt3_txphdlyreset_i
        .gt3_txphinit_in                (gt3_txphinit_i), // input wire gt3_txphinit_i
        .gt3_txphinitdone_out           (gt3_txphinitdone_i), // output wire gt3_txphinitdone_i
        //-------------------- Transmit Ports - TX Buffer Ports --------------------
        .gt3_txbufstatus_out            (gt3_txbufstatus_out), // output wire [1:0] gt3_txbufstatus_out
        //------------- Transmit Ports - TX Configurable Driver Ports --------------
        .gt3_txdiffctrl_in              (gt3_txdiffctrl_in), // input wire [3:0] gt3_txdiffctrl_in
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .gt3_txdata_in                  (gt3_txdata_in), // input wire [19:0] gt3_txdata_in
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .gt3_gtxtxn_out                 (gt3_gtxtxn_out), // output wire gt3_gtxtxn_out
        .gt3_gtxtxp_out                 (gt3_gtxtxp_out), // output wire gt3_gtxtxp_out
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .gt3_txoutclk_out               (gt3_txoutclk_i), // output wire gt3_txoutclk_i
        .gt3_txoutclkfabric_out         (gt3_txoutclkfabric_out), // output wire gt3_txoutclkfabric_out
        .gt3_txoutclkpcs_out            (gt3_txoutclkpcs_out), // output wire gt3_txoutclkpcs_out
        .gt3_txratedone_out             (gt3_txratedone_out), // output wire gt3_txratedone_out
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .gt3_txpcsreset_in              (gt3_txpcsreset_in), // input wire gt3_txpcsreset_in
        .gt3_txpmareset_in              (gt3_txpmareset_in), // input wire gt3_txpmareset_in
        .gt3_txresetdone_out            (gt3_txresetdone_i), // output wire gt3_txresetdone_i




    //____________________________COMMON PORTS________________________________
        .gt0_qplloutclk_in              (gt0_qplloutclk_in),
        .gt0_qplloutrefclk_in           (gt0_qplloutrefclk_in)

    );

assign  gt0_rxpcsreset_i                     =  tied_to_ground_i;
assign  gt0_txpcsreset_i                     =  tied_to_ground_i;
assign  gt1_rxpcsreset_i                     =  tied_to_ground_i;
assign  gt1_txpcsreset_i                     =  tied_to_ground_i;
assign  gt2_rxpcsreset_i                     =  tied_to_ground_i;
assign  gt2_txpcsreset_i                     =  tied_to_ground_i;
assign  gt3_rxpcsreset_i                     =  tied_to_ground_i;
assign  gt3_txpcsreset_i                     =  tied_to_ground_i;

    assign  gt0_rxdfelpmreset_i                  =  tied_to_ground_i;
assign  gt0_txpmareset_i                     =  tied_to_ground_i;
    assign  gt1_rxdfelpmreset_i                  =  tied_to_ground_i;
assign  gt1_txpmareset_i                     =  tied_to_ground_i;
    assign  gt2_rxdfelpmreset_i                  =  tied_to_ground_i;
assign  gt2_txpmareset_i                     =  tied_to_ground_i;
    assign  gt3_rxdfelpmreset_i                  =  tied_to_ground_i;
assign  gt3_txpmareset_i                     =  tied_to_ground_i;

assign  gt0_txsysclksel_i                    =  2'b11;
assign  gt1_txsysclksel_i                    =  2'b11;
assign  gt2_txsysclksel_i                    =  2'b11;
assign  gt3_txsysclksel_i                    =  2'b11;

assign  gt0_txresetdone_out                  =  gt0_txresetdone_i;
assign  gt0_rxresetdone_out                  =  gt0_rxresetdone_i;
assign  gt0_rxoutclk_out                     =  gt0_rxoutclk_i;
assign  gt0_txoutclk_out                     =  gt0_txoutclk_i;
assign  gt1_txresetdone_out                  =  gt1_txresetdone_i;
assign  gt1_rxresetdone_out                  =  gt1_rxresetdone_i;
assign  gt1_rxoutclk_out                     =  gt1_rxoutclk_i;
assign  gt1_txoutclk_out                     =  gt1_txoutclk_i;
assign  gt2_txresetdone_out                  =  gt2_txresetdone_i;
assign  gt2_rxresetdone_out                  =  gt2_rxresetdone_i;
assign  gt2_rxoutclk_out                     =  gt2_rxoutclk_i;
assign  gt2_txoutclk_out                     =  gt2_txoutclk_i;
assign  gt3_txresetdone_out                  =  gt3_txresetdone_i;
assign  gt3_rxresetdone_out                  =  gt3_rxresetdone_i;
assign  gt3_rxoutclk_out                     =  gt3_rxoutclk_i;
assign  gt3_txoutclk_out                     =  gt3_txoutclk_i;
assign  gt0_qpllreset_out                    =  gt0_qpllreset_t;

generate
if (EXAMPLE_USE_CHIPSCOPE == 1) 
begin : chipscope
assign  gt0_gttxreset_i                      =  gt0_gttxreset_in || gt0_gttxreset_t;
assign  gt0_gtrxreset_i                      =  gt0_gtrxreset_in || gt0_gtrxreset_t;
assign  gt0_txuserrdy_i                      =  gt0_txuserrdy_in || gt0_txuserrdy_t;
assign  gt0_rxuserrdy_i                      =  gt0_rxuserrdy_in || gt0_rxuserrdy_t;
assign  gt1_gttxreset_i                      =  gt1_gttxreset_in || gt1_gttxreset_t;
assign  gt1_gtrxreset_i                      =  gt1_gtrxreset_in || gt1_gtrxreset_t;
assign  gt1_txuserrdy_i                      =  gt1_txuserrdy_in || gt1_txuserrdy_t;
assign  gt1_rxuserrdy_i                      =  gt1_rxuserrdy_in || gt1_rxuserrdy_t;
assign  gt2_gttxreset_i                      =  gt2_gttxreset_in || gt2_gttxreset_t;
assign  gt2_gtrxreset_i                      =  gt2_gtrxreset_in || gt2_gtrxreset_t;
assign  gt2_txuserrdy_i                      =  gt2_txuserrdy_in || gt2_txuserrdy_t;
assign  gt2_rxuserrdy_i                      =  gt2_rxuserrdy_in || gt2_rxuserrdy_t;
assign  gt3_gttxreset_i                      =  gt3_gttxreset_in || gt3_gttxreset_t;
assign  gt3_gtrxreset_i                      =  gt3_gtrxreset_in || gt3_gtrxreset_t;
assign  gt3_txuserrdy_i                      =  gt3_txuserrdy_in || gt3_txuserrdy_t;
assign  gt3_rxuserrdy_i                      =  gt3_rxuserrdy_in || gt3_rxuserrdy_t;
end
endgenerate 

generate
if (EXAMPLE_USE_CHIPSCOPE == 0) 
begin : no_chipscope
assign  gt0_gttxreset_i                      =  gt0_gttxreset_t;
assign  gt0_gtrxreset_i                      =  gt0_gtrxreset_t;
assign  gt0_txuserrdy_i                      =  gt0_txuserrdy_t;
assign  gt0_rxuserrdy_i                      =  gt0_rxuserrdy_t;
assign  gt1_gttxreset_i                      =  gt1_gttxreset_t;
assign  gt1_gtrxreset_i                      =  gt1_gtrxreset_t;
assign  gt1_txuserrdy_i                      =  gt1_txuserrdy_t;
assign  gt1_rxuserrdy_i                      =  gt1_rxuserrdy_t;
assign  gt2_gttxreset_i                      =  gt2_gttxreset_t;
assign  gt2_gtrxreset_i                      =  gt2_gtrxreset_t;
assign  gt2_txuserrdy_i                      =  gt2_txuserrdy_t;
assign  gt2_rxuserrdy_i                      =  gt2_rxuserrdy_t;
assign  gt3_gttxreset_i                      =  gt3_gttxreset_t;
assign  gt3_gtrxreset_i                      =  gt3_gtrxreset_t;
assign  gt3_txuserrdy_i                      =  gt3_txuserrdy_t;
assign  gt3_rxuserrdy_i                      =  gt3_rxuserrdy_t;
end
endgenerate 


gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("TRUE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt0_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt0_txusrclk_in),
        .SOFT_RESET                     (soft_reset_tx_in),
        .QPLLREFCLKLOST                 (gt0_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt0_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt0_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt0_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (gt0_qpllreset_t),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt0_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt0_txuserrdy_t),
        .RUN_PHALIGNMENT                (gt0_run_tx_phalignment_i),
        .RESET_PHALIGNMENT              (gt0_rst_tx_phalignment_i),
        .PHALIGNMENT_DONE               (gt0_tx_phalignment_done_i),
        .RETRY_COUNTER                  ()
           );


gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("TRUE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt1_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt1_txusrclk_in),
        .SOFT_RESET                     (soft_reset_tx_in),
        .QPLLREFCLKLOST                 (gt0_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt0_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt1_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt1_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt1_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt1_txuserrdy_t),
        .RUN_PHALIGNMENT                (gt1_run_tx_phalignment_i),
        .RESET_PHALIGNMENT              (gt1_rst_tx_phalignment_i),
        .PHALIGNMENT_DONE               (gt0_tx_phalignment_done_i),
        .RETRY_COUNTER                  ()
           );


gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("TRUE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt2_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt2_txusrclk_in),
        .SOFT_RESET                     (soft_reset_tx_in),
        .QPLLREFCLKLOST                 (gt0_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt0_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt2_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt2_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt2_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt2_txuserrdy_t),
        .RUN_PHALIGNMENT                (gt2_run_tx_phalignment_i),
        .RESET_PHALIGNMENT              (gt2_rst_tx_phalignment_i),
        .PHALIGNMENT_DONE               (gt0_tx_phalignment_done_i),
        .RETRY_COUNTER                  ()
           );


gtwizard_0_TX_STARTUP_FSM #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                        // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                        // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("TRUE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt3_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (sysclk_in),
        .TXUSERCLK                      (gt3_txusrclk_in),
        .SOFT_RESET                     (soft_reset_tx_in),
        .QPLLREFCLKLOST                 (gt0_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt0_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .TXRESETDONE                    (gt3_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt3_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .TX_FSM_RESET_DONE              (gt3_tx_fsm_reset_done_out),
        .TXUSERRDY                      (gt3_txuserrdy_t),
        .RUN_PHALIGNMENT                (gt3_run_tx_phalignment_i),
        .RESET_PHALIGNMENT              (gt3_rst_tx_phalignment_i),
        .PHALIGNMENT_DONE               (gt0_tx_phalignment_done_i),
        .RETRY_COUNTER                  ()
           );





gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("TRUE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt0_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt0_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_rx_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt0_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt0_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt0_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt0_data_valid_in),
        .TXUSERRDY                      (tied_to_vcc_i),
        .GTRXRESET                      (gt0_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt0_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt0_rxuserrdy_t),
        .RUN_PHALIGNMENT                (gt0_run_rx_phalignment_i),
        .RESET_PHALIGNMENT              (gt0_rst_rx_phalignment_i),
        .PHALIGNMENT_DONE               (gt0_rx_phalignment_done_i),
        .RXDFEAGCHOLD                   (gt0_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt0_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt0_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt0_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("TRUE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt1_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt1_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_rx_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt0_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt0_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt1_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt1_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt1_data_valid_in),
        .TXUSERRDY                      (tied_to_vcc_i),
        .GTRXRESET                      (gt1_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt1_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt1_rxuserrdy_t),
        .RUN_PHALIGNMENT                (gt1_run_rx_phalignment_i),
        .RESET_PHALIGNMENT              (gt1_rst_rx_phalignment_i),
        .PHALIGNMENT_DONE               (gt0_rx_phalignment_done_i),
        .RXDFEAGCHOLD                   (gt1_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt1_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt1_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt1_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("TRUE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt2_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt2_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_rx_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt0_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt0_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt2_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt2_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt2_data_valid_in),
        .TXUSERRDY                      (tied_to_vcc_i),
        .GTRXRESET                      (gt2_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt2_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt2_rxuserrdy_t),
        .RUN_PHALIGNMENT                (gt2_run_rx_phalignment_i),
        .RESET_PHALIGNMENT              (gt2_rst_rx_phalignment_i),
        .PHALIGNMENT_DONE               (gt0_rx_phalignment_done_i),
        .RXDFEAGCHOLD                   (gt2_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt2_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt2_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt2_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

gtwizard_0_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("TRUE"),                           // the TX and RX Reset FSMs must 
           .RX_QPLL_USED             ("TRUE"),                           // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("TRUE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt3_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (sysclk_in),
        .RXUSERCLK                      (gt3_rxusrclk_in),
        .SOFT_RESET                     (soft_reset_rx_in),
        .DONT_RESET_ON_DATA_ERROR       (dont_reset_on_data_error_in),
        .QPLLREFCLKLOST                 (gt0_qpllrefclklost_in),
        .CPLLREFCLKLOST                 (tied_to_ground_i),
        .QPLLLOCK                       (gt0_qplllock_in),
        .CPLLLOCK                       (tied_to_vcc_i),
        .RXRESETDONE                    (gt3_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt3_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (gt3_data_valid_in),
        .TXUSERRDY                      (tied_to_vcc_i),
        .GTRXRESET                      (gt3_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (gt3_rx_fsm_reset_done_out),
        .RXUSERRDY                      (gt3_rxuserrdy_t),
        .RUN_PHALIGNMENT                (gt3_run_rx_phalignment_i),
        .RESET_PHALIGNMENT              (gt3_rst_rx_phalignment_i),
        .PHALIGNMENT_DONE               (gt0_rx_phalignment_done_i),
        .RXDFEAGCHOLD                   (gt3_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt3_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt3_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt3_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

  always @(posedge sysclk_in)
  begin
        if(gt0_gtrxreset_i)
        begin
          gt0_rx_cdrlocked       <= `DLY    1'b0;
          gt0_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt0_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt0_rx_cdrlocked       <= `DLY    1'b1;
          gt0_rx_cdrlock_counter <= `DLY    gt0_rx_cdrlock_counter;
        end
        else
          gt0_rx_cdrlock_counter <= `DLY    gt0_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt1_gtrxreset_i)
        begin
          gt1_rx_cdrlocked       <= `DLY    1'b0;
          gt1_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt1_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt1_rx_cdrlocked       <= `DLY    1'b1;
          gt1_rx_cdrlock_counter <= `DLY    gt1_rx_cdrlock_counter;
        end
        else
          gt1_rx_cdrlock_counter <= `DLY    gt1_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt2_gtrxreset_i)
        begin
          gt2_rx_cdrlocked       <= `DLY    1'b0;
          gt2_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt2_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt2_rx_cdrlocked       <= `DLY    1'b1;
          gt2_rx_cdrlock_counter <= `DLY    gt2_rx_cdrlock_counter;
        end
        else
          gt2_rx_cdrlock_counter <= `DLY    gt2_rx_cdrlock_counter + 1;
  end 

  always @(posedge sysclk_in)
  begin
        if(gt3_gtrxreset_i)
        begin
          gt3_rx_cdrlocked       <= `DLY    1'b0;
          gt3_rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (gt3_rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          gt3_rx_cdrlocked       <= `DLY    1'b1;
          gt3_rx_cdrlock_counter <= `DLY    gt3_rx_cdrlock_counter;
        end
        else
          gt3_rx_cdrlock_counter <= `DLY    gt3_rx_cdrlock_counter + 1;
  end 

assign  gt0_recclk_stable_i                  =  gt0_rx_cdrlocked;
assign  gt1_recclk_stable_i                  =  gt1_rx_cdrlocked;
assign  gt2_recclk_stable_i                  =  gt2_rx_cdrlocked;
assign  gt3_recclk_stable_i                  =  gt3_rx_cdrlocked;



//   --------------------------- TX Buffer Bypass Logic --------------------
//   The TX SYNC Module drives the ports needed to Bypass the TX Buffer.
//   Include the TX SYNC module in your own design if TX Buffer is bypassed.

//Manual
   gtwizard_0_TX_MANUAL_PHASE_ALIGN #
   (
     .NUMBER_OF_LANES	  (4),
     .MASTER_LANE_ID      (0)
   )
   gt0_tx_manual_phase_i 
   (
        .STABLE_CLOCK                   (sysclk_in),
        .RESET_PHALIGNMENT              (U0_rst_tx_phalignment_i),   
        .RUN_PHALIGNMENT                (U0_run_tx_phalignment_i),      
        .PHASE_ALIGNMENT_DONE           (gt0_tx_phalignment_done_i),
        .TXDLYSRESET                    (U0_TXDLYSRESET),
        .TXDLYSRESETDONE                (U0_TXDLYSRESETDONE),
        .TXPHINIT                       (U0_TXPHINIT),
        .TXPHINITDONE                   (U0_TXPHINITDONE),
        .TXPHALIGN                      (U0_TXPHALIGN),
        .TXPHALIGNDONE                  (U0_TXPHALIGNDONE),
        .TXDLYEN                        (U0_TXDLYEN)
   );

assign  gt0_txphdlyreset_i                   =  tied_to_ground_i;
assign  gt0_txphalignen_i                    =  tied_to_vcc_i;
assign  gt0_txdlysreset_i                    =  U0_TXDLYSRESET[0];
assign  gt0_txphinit_i                       =  U0_TXPHINIT[0];
assign  gt0_txphalign_i                      =  U0_TXPHALIGN[0];
assign  gt0_txdlyen_i                        =  U0_TXDLYEN[0];
assign  U0_TXDLYSRESETDONE[0]                =  gt0_txdlysresetdone_i;
assign  U0_TXPHINITDONE[0]                   =  gt0_txphinitdone_i;
assign  U0_TXPHALIGNDONE[0]                  =  gt0_txphaligndone_i;



 
assign  gt1_txdlysreset_i                    =  U0_TXDLYSRESET[1];
assign  gt1_txphinit_i                       =  U0_TXPHINIT[1];
assign  gt1_txphalign_i                      =  U0_TXPHALIGN[1];
assign  gt1_txphalignen_i                    =  tied_to_vcc_i;
assign  gt1_txphdlyreset_i                   =  tied_to_ground_i;
assign  gt1_txdlyen_i                        =  tied_to_ground_i;
assign  U0_TXDLYSRESETDONE[1]                =  gt1_txdlysresetdone_i;
assign  U0_TXPHINITDONE[1]                   =  gt1_txphinitdone_i;
assign  U0_TXPHALIGNDONE[1]                  =  gt1_txphaligndone_i;


 
assign  gt2_txdlysreset_i                    =  U0_TXDLYSRESET[2];
assign  gt2_txphinit_i                       =  U0_TXPHINIT[2];
assign  gt2_txphalign_i                      =  U0_TXPHALIGN[2];
assign  gt2_txphalignen_i                    =  tied_to_vcc_i;
assign  gt2_txphdlyreset_i                   =  tied_to_ground_i;
assign  gt2_txdlyen_i                        =  tied_to_ground_i;
assign  U0_TXDLYSRESETDONE[2]                =  gt2_txdlysresetdone_i;
assign  U0_TXPHINITDONE[2]                   =  gt2_txphinitdone_i;
assign  U0_TXPHALIGNDONE[2]                  =  gt2_txphaligndone_i;


 
assign  gt3_txdlysreset_i                    =  U0_TXDLYSRESET[3];
assign  gt3_txphinit_i                       =  U0_TXPHINIT[3];
assign  gt3_txphalign_i                      =  U0_TXPHALIGN[3];
assign  gt3_txphalignen_i                    =  tied_to_vcc_i;
assign  gt3_txphdlyreset_i                   =  tied_to_ground_i;
assign  gt3_txdlyen_i                        =  tied_to_ground_i;
assign  U0_TXDLYSRESETDONE[3]                =  gt3_txdlysresetdone_i;
assign  U0_TXPHINITDONE[3]                   =  gt3_txphinitdone_i;
assign  U0_TXPHALIGNDONE[3]                  =  gt3_txphaligndone_i;



  assign  U0_run_tx_phalignment_i    =  gt0_run_tx_phalignment_i 
 
                                             && gt1_run_tx_phalignment_i
 
                                             && gt2_run_tx_phalignment_i
 
                                             && gt3_run_tx_phalignment_i
                                             ;

    assign U0_rst_tx_phalignment_i   =  gt0_rst_tx_phalignment_i 
 
                                             || gt1_rst_tx_phalignment_i
 
                                             || gt2_rst_tx_phalignment_i
 
                                             || gt3_rst_tx_phalignment_i
                                             ;




//   --------------------------- RX Buffer Bypass Logic --------------------
//   The RX SYNC Module drives the ports needed to Bypass the RX Buffer.
//   Include the RX SYNC module in your own design if RX Buffer is bypassed.

//Manual
   gtwizard_0_RX_MANUAL_PHASE_ALIGN #
   (
     .NUMBER_OF_LANES	  (4),
     .MASTER_LANE_ID      (0)
   )
   gt0_rx_manual_phase_i 
   (
        .STABLE_CLOCK                   (sysclk_in),
        .RESET_PHALIGNMENT              (U0_rst_rx_phalignment_i),   
        .RUN_PHALIGNMENT                (U0_run_rx_phalignment_i),      
        .PHASE_ALIGNMENT_DONE           (gt0_rx_phalignment_done_i),
        .RXDLYSRESET                    (U0_RXDLYSRESET),
        .RXDLYSRESETDONE                (U0_RXDLYSRESETDONE),
        .RXPHALIGN                      (U0_RXPHALIGN),
        .RXPHALIGNDONE                  (U0_RXPHALIGNDONE),
        .RXDLYEN                        (U0_RXDLYEN)
   );

assign  gt0_rxphdlyreset_i                   =  tied_to_ground_i;
assign  gt0_rxphalignen_i                    =  tied_to_vcc_i;
assign  gt0_rxdlysreset_i                    =  U0_RXDLYSRESET[0];
assign  gt0_rxphalign_i                      =  U0_RXPHALIGN[0];
assign  gt0_rxdlyen_i                        =  U0_RXDLYEN[0];
assign  U0_RXDLYSRESETDONE[0]                =  gt0_rxdlysresetdone_i;
assign  U0_RXPHALIGNDONE[0]                  =  gt0_rxphaligndone_i;



 
assign  gt1_rxdlysreset_i                    =  U0_RXDLYSRESET[1];
assign  gt1_rxphalign_i                      =  U0_RXPHALIGN[1];
assign  gt1_rxphalignen_i                    =  tied_to_vcc_i;
assign  gt1_rxphdlyreset_i                   =  tied_to_ground_i;
assign  gt1_rxdlyen_i                        =  tied_to_ground_i;
assign  U0_RXDLYSRESETDONE[1]                =  gt1_rxdlysresetdone_i;
assign  U0_RXPHALIGNDONE[1]                  =  gt1_rxphaligndone_i;


 
assign  gt2_rxdlysreset_i                    =  U0_RXDLYSRESET[2];
assign  gt2_rxphalign_i                      =  U0_RXPHALIGN[2];
assign  gt2_rxphalignen_i                    =  tied_to_vcc_i;
assign  gt2_rxphdlyreset_i                   =  tied_to_ground_i;
assign  gt2_rxdlyen_i                        =  tied_to_ground_i;
assign  U0_RXDLYSRESETDONE[2]                =  gt2_rxdlysresetdone_i;
assign  U0_RXPHALIGNDONE[2]                  =  gt2_rxphaligndone_i;


 
assign  gt3_rxdlysreset_i                    =  U0_RXDLYSRESET[3];
assign  gt3_rxphalign_i                      =  U0_RXPHALIGN[3];
assign  gt3_rxphalignen_i                    =  tied_to_vcc_i;
assign  gt3_rxphdlyreset_i                   =  tied_to_ground_i;
assign  gt3_rxdlyen_i                        =  tied_to_ground_i;
assign  U0_RXDLYSRESETDONE[3]                =  gt3_rxdlysresetdone_i;
assign  U0_RXPHALIGNDONE[3]                  =  gt3_rxphaligndone_i;



  assign  U0_run_rx_phalignment_i    =  gt0_run_rx_phalignment_i 
 
                                             && gt1_run_rx_phalignment_i
 
                                             && gt2_run_rx_phalignment_i
 
                                             && gt3_run_rx_phalignment_i
                                             ;

    assign U0_rst_rx_phalignment_i    =  gt0_rst_rx_phalignment_i 
 
                                             || gt1_rst_rx_phalignment_i
 
                                             || gt2_rst_rx_phalignment_i
 
                                             || gt3_rst_rx_phalignment_i
                                             ;


endmodule


